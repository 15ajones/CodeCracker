
module CodeCracker (
	accelerometer_spi_0_external_interface_I2C_SDAT,
	accelerometer_spi_0_external_interface_I2C_SCLK,
	accelerometer_spi_0_external_interface_G_SENSOR_CS_N,
	accelerometer_spi_0_external_interface_G_SENSOR_INT,
	button_external_connection_export,
	clk_clk,
	hex0_external_connection_export,
	hex1_external_connection_export,
	hex2_external_connection_export,
	hex3_external_connection_export,
	hex4_external_connection_export,
	hex5_external_connection_export,
	led_external_connection_export,
	reset_reset_n,
	switch_external_connection_export,
	uart_0_external_connection_rxd,
	uart_0_external_connection_txd);	

	inout		accelerometer_spi_0_external_interface_I2C_SDAT;
	output		accelerometer_spi_0_external_interface_I2C_SCLK;
	output		accelerometer_spi_0_external_interface_G_SENSOR_CS_N;
	input		accelerometer_spi_0_external_interface_G_SENSOR_INT;
	input	[3:0]	button_external_connection_export;
	input		clk_clk;
	output	[6:0]	hex0_external_connection_export;
	output	[6:0]	hex1_external_connection_export;
	output	[6:0]	hex2_external_connection_export;
	output	[6:0]	hex3_external_connection_export;
	output	[6:0]	hex4_external_connection_export;
	output	[6:0]	hex5_external_connection_export;
	output	[9:0]	led_external_connection_export;
	input		reset_reset_n;
	input	[9:0]	switch_external_connection_export;
	input		uart_0_external_connection_rxd;
	output		uart_0_external_connection_txd;
endmodule
